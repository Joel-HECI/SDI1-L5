-- (110) Realizar la operación XOR de X, Y y D
