-- (101) Realizar la operación OR de los dos números X y Y
